// 简单的testbench，观测寄存器链传递
`timescale 1ns/1ps
module tb;
    reg clk;
    reg resetn;
    reg  [7:0] switch;
    wire [15:0] led;

    initial begin
        clk = 1'b0;
        resetn = 1'b0;
        #2000;
        resetn = 1'b1;
    end
    always #5 clk = ~clk;

    initial begin
        // 可自定义测试输入
        switch = ~(8'h5);
    end

    soc_mini_top dut (
        .resetn (resetn),
        .clk    (clk),
        .led    (led),
        .switch (switch)
    );

    initial begin
        $monitor($time, " led = %h", led);
        #5000;
        $finish;
    end
endmodule
